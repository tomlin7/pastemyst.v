module tests

