module types

pub struct RawTime {
	result int [json: result]
}