module pastemyst

import src
import tests


import json
import net.http

const main_endpoint  = "https://paste.myst.rs/api/v2"
