module pastemyst

import src
import tests