module types

pub struct RawTime {
pub:
	result int [json: result]
}