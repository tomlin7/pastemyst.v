module pastemyst

/**
 * The base endpoint to make requests to.
 */
pub const main_endpoint  = "https://paste.myst.rs/api/v2"
