module types

/**
 * Represents an timestamp conversion result.
 *
 * @see https://paste.myst.rs/api-docs/objects
 */
pub struct RawTime {
pub:
	/**
	 * The result of the conversion.
	 */
	result int [json: result]
}