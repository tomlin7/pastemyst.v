module pastemyst

pub const main_endpoint  = "https://paste.myst.rs/api/v2"
