module pastemyst