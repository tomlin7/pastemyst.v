module tests

import { data } from "./pastemyst";

fn test_hello() {
    assert hello() == 'Hello world'
}


