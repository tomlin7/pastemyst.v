module types

import json

pub struct RawTime {
	result int [json: result]
}