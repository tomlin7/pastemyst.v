module pastemyst

// tests

// get public paste
// println("Getting paste")
// println(get_paste(id: '99is6n23'))

// get private paste
// println("Getting private paste")
// println(get_paste(id: 'xc9mvyaq', token: 'token'))

// create public paste 

// fn main () {
//     mut new_pasty := Pasty {
//         language: "autodetect"
//         title   : "test"
//         code    : "print('test')"
//     }
//     mut new_paste := Paste {
//         title   : "test"
//         pasties : [new_pasty]
//     }

//     mut result := create_paste(paste: new_paste) ?
//     print(result.str())
// }

// create private paste 

// fn main () {
//     mut new_pasty := Pasty {
//         language: "autodetect"
//         title   : "test"
//         code    : "print('test')"
//     }
//     mut new_paste := Paste {
//         title   : "test"
//         pasties : [new_pasty]
//     }

//     mut result := create_paste(paste: new_paste, token: "token") ?
//     print(result.str())
// }

// delete a paste

