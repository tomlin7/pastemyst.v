module pastemyst

// import types
// import endpoints 

// import tests


import json
import net.http

pub const main_endpoint  = "https://paste.myst.rs/api/v2"
