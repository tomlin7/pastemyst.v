module pastemyst

// import types
// import endpoints 

// import tests

pub const main_endpoint  = "https://paste.myst.rs/api/v2"
