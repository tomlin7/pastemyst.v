module pastemyst

import src