module tests